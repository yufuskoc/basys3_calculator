`timescale 1ns / 1ps

module prime(clk, reset, number, result);

input clk;
input reset;
input [8:0]number;
output reg result;
  
always @(posedge clk) begin
    if(number==0)result=0;
    else if(number==1)result=0;
    else if(number==2)result=1;
    else if(number==3)result=1;
    else if(number==4)result=0;
    else if(number==5)result=1;
    else if(number==6)result=0;
    else if(number==7)result=1;
    else if(number==8)result=0;
    else if(number==9)result=0;
    else if(number==10)result=0;
    else if(number==11)result=1;
    else if(number==12)result=0;
    else if(number==13)result=1;
    else if(number==14)result=0;
    else if(number==15)result=0;
    else if(number==16)result=0;
    else if(number==17)result=1;
    else if(number==18)result=0;
    else if(number==19)result=1;
    else if(number==20)result=0;
    else if(number==21)result=0;
    else if(number==22)result=0;
    else if(number==23)result=1;
    else if(number==24)result=0;
    else if(number==25)result=0;
    else if(number==26)result=0;
    else if(number==27)result=0;
    else if(number==28)result=0;
    else if(number==29)result=1;
    else if(number==30)result=0;
    else if(number==31)result=1;
    else if(number==32)result=0;
    else if(number==33)result=0;
    else if(number==34)result=0;
    else if(number==35)result=0;
    else if(number==36)result=0;
    else if(number==37)result=1;
    else if(number==38)result=0;
    else if(number==39)result=0;
    else if(number==40)result=0;
    else if(number==41)result=1;
    else if(number==42)result=0;
    else if(number==43)result=1;
    else if(number==44)result=0;
    else if(number==45)result=0;
    else if(number==46)result=0;
    else if(number==47)result=1;
    else if(number==48)result=0;
    else if(number==49)result=0;
    else if(number==50)result=0;
    else if(number==51)result=0;
    else if(number==52)result=0;
    else if(number==53)result=1;
    else if(number==54)result=0;
    else if(number==55)result=0;
    else if(number==56)result=0;
    else if(number==57)result=0;
    else if(number==58)result=0;
    else if(number==59)result=1;
    else if(number==60)result=0;
    else if(number==61)result=1;
    else if(number==62)result=0;
    else if(number==63)result=0;
    else if(number==64)result=0;
    else if(number==65)result=0;
    else if(number==66)result=0;
    else if(number==67)result=1;
    else if(number==68)result=0;
    else if(number==69)result=0;
    else if(number==70)result=0;
    else if(number==71)result=1;
    else if(number==72)result=0;
    else if(number==73)result=1;
    else if(number==74)result=0;
    else if(number==75)result=0;
    else if(number==76)result=0;
    else if(number==77)result=0;
    else if(number==78)result=0;
    else if(number==79)result=1;
    else if(number==80)result=0;
    else if(number==81)result=0;
    else if(number==82)result=0;
    else if(number==83)result=1;
    else if(number==84)result=0;
    else if(number==85)result=0;
    else if(number==86)result=0;
    else if(number==87)result=0;
    else if(number==88)result=0;
    else if(number==89)result=1;
    else if(number==90)result=0;
    else if(number==91)result=0;
    else if(number==92)result=0;
    else if(number==93)result=0;
    else if(number==94)result=0;
    else if(number==95)result=0;
    else if(number==96)result=0;
    else if(number==97)result=1;
    else if(number==98)result=0;
    else if(number==99)result=0;
    else if(number==100)result=0;
    else if(number==101)result=1;
    else if(number==102)result=0;
    else if(number==103)result=1;
    else if(number==104)result=0;
    else if(number==105)result=0;
    else if(number==106)result=0;
    else if(number==107)result=1;
    else if(number==108)result=0;
    else if(number==109)result=1;
    else if(number==110)result=0;
    else if(number==111)result=0;
    else if(number==112)result=0;
    else if(number==113)result=1;
    else if(number==114)result=0;
    else if(number==115)result=0;
    else if(number==116)result=0;
    else if(number==117)result=0;
    else if(number==118)result=0;
    else if(number==119)result=0;
    else if(number==120)result=0;
    else if(number==121)result=0;
    else if(number==122)result=0;
    else if(number==123)result=0;
    else if(number==124)result=0;
    else if(number==125)result=0;
    else if(number==126)result=0;
    else if(number==127)result=1;
    else if(number==128)result=0;
    else if(number==129)result=0;
    else if(number==130)result=0;
    else if(number==131)result=1;
    else if(number==132)result=0;
    else if(number==133)result=0;
    else if(number==134)result=0;
    else if(number==135)result=0;
    else if(number==136)result=0;
    else if(number==137)result=1;
    else if(number==138)result=0;
    else if(number==139)result=1;
    else if(number==140)result=0;
    else if(number==141)result=0;
    else if(number==142)result=0;
    else if(number==143)result=0;
    else if(number==144)result=0;
    else if(number==145)result=0;
    else if(number==146)result=0;
    else if(number==147)result=0;
    else if(number==148)result=0;
    else if(number==149)result=1;
    else if(number==150)result=0;
    else if(number==151)result=1;
    else if(number==152)result=0;
    else if(number==153)result=0;
    else if(number==154)result=0;
    else if(number==155)result=0;
    else if(number==156)result=0;
    else if(number==157)result=1;
    else if(number==158)result=0;
    else if(number==159)result=0;
    else if(number==160)result=0;
    else if(number==161)result=0;
    else if(number==162)result=0;
    else if(number==163)result=1;
    else if(number==164)result=0;
    else if(number==165)result=0;
    else if(number==166)result=0;
    else if(number==167)result=1;
    else if(number==168)result=0;
    else if(number==169)result=0;
    else if(number==170)result=0;
    else if(number==171)result=0;
    else if(number==172)result=0;
    else if(number==173)result=1;
    else if(number==174)result=0;
    else if(number==175)result=0;
    else if(number==176)result=0;
    else if(number==177)result=0;
    else if(number==178)result=0;
    else if(number==179)result=1;
    else if(number==180)result=0;
    else if(number==181)result=1;
    else if(number==182)result=0;
    else if(number==183)result=0;
    else if(number==184)result=0;
    else if(number==185)result=0;
    else if(number==186)result=0;
    else if(number==187)result=0;
    else if(number==188)result=0;
    else if(number==189)result=0;
    else if(number==190)result=0;
    else if(number==191)result=1;
    else if(number==192)result=0;
    else if(number==193)result=1;
    else if(number==194)result=0;
    else if(number==195)result=0;
    else if(number==196)result=0;
    else if(number==197)result=1;
    else if(number==198)result=0;
    else if(number==199)result=1;
    else if(number==200)result=0;
    else if(number==201)result=0;
    else if(number==202)result=0;
    else if(number==203)result=0;
    else if(number==204)result=0;
    else if(number==205)result=0;
    else if(number==206)result=0;
    else if(number==207)result=0;
    else if(number==208)result=0;
    else if(number==209)result=0;
    else if(number==210)result=0;
    else if(number==211)result=1;
    else if(number==212)result=0;
    else if(number==213)result=0;
    else if(number==214)result=0;
    else if(number==215)result=0;
    else if(number==216)result=0;
    else if(number==217)result=0;
    else if(number==218)result=0;
    else if(number==219)result=0;
    else if(number==220)result=0;
    else if(number==221)result=0;
    else if(number==222)result=0;
    else if(number==223)result=1;
    else if(number==224)result=0;
    else if(number==225)result=0;
    else if(number==226)result=0;
    else if(number==227)result=1;
    else if(number==228)result=0;
    else if(number==229)result=1;
    else if(number==230)result=0;
    else if(number==231)result=0;
    else if(number==232)result=0;
    else if(number==233)result=1;
    else if(number==234)result=0;
    else if(number==235)result=0;
    else if(number==236)result=0;
    else if(number==237)result=0;
    else if(number==238)result=0;
    else if(number==239)result=1;
    else if(number==240)result=0;
    else if(number==241)result=1;
    else if(number==242)result=0;
    else if(number==243)result=0;
    else if(number==244)result=0;
    else if(number==245)result=0;
    else if(number==246)result=0;
    else if(number==247)result=0;
    else if(number==248)result=0;
    else if(number==249)result=0;
    else if(number==250)result=0;
    else if(number==251)result=1;
    else if(number==252)result=0;
    else if(number==253)result=0;
    else if(number==254)result=0;
    else if(number==255)result=0;
    else if(number==256)result=0;
    else if(number==257)result=1;
    else if(number==258)result=0;
    else if(number==259)result=0;
    else if(number==260)result=0;
    else if(number==261)result=0;
    else if(number==262)result=0;
    else if(number==263)result=1;
    else if(number==264)result=0;
    else if(number==265)result=0;
    else if(number==266)result=0;
    else if(number==267)result=0;
    else if(number==268)result=0;
    else if(number==269)result=1;
    else if(number==270)result=0;
    else if(number==271)result=1;
    else if(number==272)result=0;
    else if(number==273)result=0;
    else if(number==274)result=0;
    else if(number==275)result=0;
    else if(number==276)result=0;
    else if(number==277)result=1;
    else if(number==278)result=0;
    else if(number==279)result=0;
    else if(number==280)result=0;
    else if(number==281)result=1;
    else if(number==282)result=0;
    else if(number==283)result=1;
    else if(number==284)result=0;
    else if(number==285)result=0;
    else if(number==286)result=0;
    else if(number==287)result=0;
    else if(number==288)result=0;
    else if(number==289)result=0;
    else if(number==290)result=0;
    else if(number==291)result=0;
    else if(number==292)result=0;
    else if(number==293)result=1;
    else if(number==294)result=0;
    else if(number==295)result=0;
    else if(number==296)result=0;
    else if(number==297)result=0;
    else if(number==298)result=0;
    else if(number==299)result=0;
    else if(number==300)result=0;
    else if(number==301)result=0;
    else if(number==302)result=0;
    else if(number==303)result=0;
    else if(number==304)result=0;
    else if(number==305)result=0;
    else if(number==306)result=0;
    else if(number==307)result=1;
    else if(number==308)result=0;
    else if(number==309)result=0;
    else if(number==310)result=0;
    else if(number==311)result=1;
    else if(number==312)result=0;
    else if(number==313)result=1;
    else if(number==314)result=0;
    else if(number==315)result=0;
    else if(number==316)result=0;
    else if(number==317)result=1;
    else if(number==318)result=0;
    else if(number==319)result=0;
    else if(number==320)result=0;
    else if(number==321)result=0;
    else if(number==322)result=0;
    else if(number==323)result=0;
    else if(number==324)result=0;
    else if(number==325)result=0;
    else if(number==326)result=0;
    else if(number==327)result=0;
    else if(number==328)result=0;
    else if(number==329)result=0;
    else if(number==330)result=0;
    else if(number==331)result=1;
    else if(number==332)result=0;
    else if(number==333)result=0;
    else if(number==334)result=0;
    else if(number==335)result=0;
    else if(number==336)result=0;
    else if(number==337)result=1;
    else if(number==338)result=0;
    else if(number==339)result=0;
    else if(number==340)result=0;
    else if(number==341)result=0;
    else if(number==342)result=0;
    else if(number==343)result=0;
    else if(number==344)result=0;
    else if(number==345)result=0;
    else if(number==346)result=0;
    else if(number==347)result=1;
    else if(number==348)result=0;
    else if(number==349)result=1;
    else if(number==350)result=0;
    else if(number==351)result=0;
    else if(number==352)result=0;
    else if(number==353)result=1;
    else if(number==354)result=0;
    else if(number==355)result=0;
    else if(number==356)result=0;
    else if(number==357)result=0;
    else if(number==358)result=0;
    else if(number==359)result=1;
    else if(number==360)result=0;
    
end

endmodule